*Model Description
.param VDD = 1.8
.param temp=27


*Including sky130 library files
.lib "sky130_fd_pr/models/sky130.lib.spice" tt


*Netlist Description


XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.15
XM2 out in 0 0 sky130_fd_pr__nfet_01v8 w=0.36 l=0.15


Cload out 0 50fF

Vdd vdd 0 {VDD}
Vin in 0 DC 0

*simulation commands

.op

* Batch-control: run DC sweep and write VTC to file
.control
  set filetype=ascii
  echo "Running inverter DC sweep for VDD={VDD}..."
  dc Vin 0 {VDD} 0.001
  wrdata vtc.dat v(in) v(out)
  quit
.endc

.end
